
module gcd ( a_in, b_in, start, reset_n, clk, result, done );
  input [31:0] a_in;
  input [31:0] b_in;
  output [31:0] result;
  input start, reset_n, clk;
  output done;
  wire   N58, N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71,
         N72, N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85,
         N86, N87, N88, N89, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, n6, n58, n59, n60, n61, n62, n63, n64, n65, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613;
  wire   [31:0] reg_a;
  wire   [31:0] reg_b;
  wire   [1:0] gcd_ns;

  DFFARX1 \reg_a_reg[0]  ( .D(N58), .CLK(clk), .RSTB(n358), .Q(reg_a[0]), .QN(
        n270) );
  DFFARX1 \reg_a_reg[29]  ( .D(N87), .CLK(clk), .RSTB(n352), .Q(reg_a[29]), 
        .QN(n198) );
  DFFARX1 \reg_a_reg[30]  ( .D(N88), .CLK(clk), .RSTB(n353), .Q(reg_a[30]), 
        .QN(n197) );
  DFFARX1 \reg_b_reg[7]  ( .D(N99), .CLK(clk), .RSTB(n356), .Q(reg_b[7]), .QN(
        n240) );
  DFFARX1 \reg_a_reg[1]  ( .D(N59), .CLK(clk), .RSTB(n357), .Q(reg_a[1]), .QN(
        n602) );
  DFFARX1 \reg_a_reg[7]  ( .D(N65), .CLK(clk), .RSTB(n356), .Q(reg_a[7]), .QN(
        n144) );
  DFFARX1 \reg_b_reg[16]  ( .D(N108), .CLK(clk), .RSTB(n346), .QN(n261) );
  DFFARX1 \reg_a_reg[3]  ( .D(N61), .CLK(clk), .RSTB(n354), .Q(reg_a[3]), .QN(
        n235) );
  DFFARX1 \gcd_ps_reg[0]  ( .D(gcd_ns[0]), .CLK(clk), .RSTB(n358), .Q(n227), 
        .QN(n67) );
  DFFARX1 \reg_b_reg[6]  ( .D(N98), .CLK(clk), .RSTB(n355), .Q(reg_b[6]), .QN(
        n230) );
  DFFARX1 \reg_b_reg[3]  ( .D(N95), .CLK(clk), .RSTB(n354), .Q(reg_b[3]), .QN(
        n178) );
  DFFARX1 \reg_b_reg[2]  ( .D(N94), .CLK(clk), .RSTB(n353), .Q(reg_b[2]), .QN(
        n219) );
  DFFARX1 \gcd_ps_reg[1]  ( .D(gcd_ns[1]), .CLK(clk), .RSTB(n356), .QN(n100)
         );
  DFFARX1 \reg_a_reg[10]  ( .D(N68), .CLK(clk), .RSTB(n343), .Q(reg_a[10]), 
        .QN(n196) );
  DFFARX1 \reg_b_reg[22]  ( .D(N114), .CLK(clk), .RSTB(n349), .Q(reg_b[22]), 
        .QN(n225) );
  DFFARX1 \reg_a_reg[16]  ( .D(N74), .CLK(clk), .RSTB(n346), .Q(reg_a[16]), 
        .QN(n216) );
  DFFARX1 \reg_a_reg[21]  ( .D(N79), .CLK(clk), .RSTB(n348), .Q(reg_a[21]), 
        .QN(n214) );
  DFFARX1 \reg_b_reg[17]  ( .D(N109), .CLK(clk), .RSTB(n346), .Q(reg_b[17]), 
        .QN(n210) );
  DFFARX1 \reg_b_reg[21]  ( .D(N113), .CLK(clk), .RSTB(n348), .Q(reg_b[21]), 
        .QN(n220) );
  DFFARX1 \reg_b_reg[8]  ( .D(N100), .CLK(clk), .RSTB(n342), .Q(reg_b[8]), 
        .QN(n212) );
  DFFARX1 \reg_b_reg[5]  ( .D(N97), .CLK(clk), .RSTB(n355), .Q(reg_b[5]), .QN(
        n215) );
  DFFARX1 \reg_a_reg[2]  ( .D(N60), .CLK(clk), .RSTB(n353), .QN(n189) );
  DFFARX1 \reg_b_reg[0]  ( .D(N92), .CLK(clk), .RSTB(n357), .Q(n176), .QN(n234) );
  DFFARX1 \reg_a_reg[5]  ( .D(N63), .CLK(clk), .RSTB(n355), .Q(reg_a[5]), .QN(
        n147) );
  DFFARX1 \result_reg[8]  ( .D(n68), .CLK(clk), .RSTB(n342), .Q(result[8]) );
  DFFARX1 \result_reg[9]  ( .D(n69), .CLK(clk), .RSTB(n342), .Q(result[9]) );
  DFFARX1 \result_reg[13]  ( .D(n73), .CLK(clk), .RSTB(n344), .Q(result[13])
         );
  DFFARX1 \result_reg[12]  ( .D(n72), .CLK(clk), .RSTB(n344), .Q(result[12])
         );
  DFFARX1 \result_reg[11]  ( .D(n71), .CLK(clk), .RSTB(n343), .Q(result[11])
         );
  DFFARX1 \result_reg[10]  ( .D(n70), .CLK(clk), .RSTB(n343), .Q(result[10])
         );
  DFFARX1 \result_reg[0]  ( .D(n99), .CLK(clk), .RSTB(n357), .Q(result[0]) );
  DFFARX1 \result_reg[31]  ( .D(n97), .CLK(clk), .RSTB(n356), .Q(result[31])
         );
  DFFARX1 \result_reg[30]  ( .D(n90), .CLK(clk), .RSTB(n353), .Q(result[30])
         );
  DFFARX1 \result_reg[29]  ( .D(n89), .CLK(clk), .RSTB(n352), .Q(result[29])
         );
  DFFARX1 \result_reg[28]  ( .D(n88), .CLK(clk), .RSTB(n352), .Q(result[28])
         );
  DFFARX1 \result_reg[27]  ( .D(n87), .CLK(clk), .RSTB(n351), .Q(result[27])
         );
  DFFARX1 \result_reg[26]  ( .D(n86), .CLK(clk), .RSTB(n351), .Q(result[26])
         );
  DFFARX1 \result_reg[25]  ( .D(n85), .CLK(clk), .RSTB(n350), .Q(result[25])
         );
  DFFARX1 \result_reg[24]  ( .D(n84), .CLK(clk), .RSTB(n350), .Q(result[24])
         );
  DFFARX1 \result_reg[23]  ( .D(n83), .CLK(clk), .RSTB(n349), .Q(result[23])
         );
  DFFARX1 \result_reg[22]  ( .D(n82), .CLK(clk), .RSTB(n349), .Q(result[22])
         );
  DFFARX1 \result_reg[21]  ( .D(n81), .CLK(clk), .RSTB(n348), .Q(result[21])
         );
  DFFARX1 \result_reg[20]  ( .D(n80), .CLK(clk), .RSTB(n348), .Q(result[20])
         );
  DFFARX1 \result_reg[19]  ( .D(n79), .CLK(clk), .RSTB(n347), .Q(result[19])
         );
  DFFARX1 \result_reg[18]  ( .D(n78), .CLK(clk), .RSTB(n347), .Q(result[18])
         );
  DFFARX1 \result_reg[17]  ( .D(n77), .CLK(clk), .RSTB(n346), .Q(result[17])
         );
  DFFARX1 \result_reg[16]  ( .D(n76), .CLK(clk), .RSTB(n346), .Q(result[16])
         );
  DFFARX1 \result_reg[15]  ( .D(n75), .CLK(clk), .RSTB(n345), .Q(result[15])
         );
  DFFARX1 \result_reg[14]  ( .D(n74), .CLK(clk), .RSTB(n345), .Q(result[14])
         );
  DFFARX1 \result_reg[7]  ( .D(n96), .CLK(clk), .RSTB(n356), .Q(result[7]) );
  DFFARX1 \result_reg[6]  ( .D(n95), .CLK(clk), .RSTB(n355), .Q(result[6]) );
  DFFARX1 \result_reg[5]  ( .D(n94), .CLK(clk), .RSTB(n355), .Q(result[5]) );
  DFFARX1 \result_reg[4]  ( .D(n93), .CLK(clk), .RSTB(n354), .Q(result[4]) );
  DFFARX1 \result_reg[3]  ( .D(n92), .CLK(clk), .RSTB(n354), .Q(result[3]) );
  DFFARX1 \result_reg[2]  ( .D(n91), .CLK(clk), .RSTB(n353), .Q(result[2]) );
  DFFARX1 \result_reg[1]  ( .D(n98), .CLK(clk), .RSTB(n357), .Q(result[1]) );
  DFFARX1 \reg_b_reg[28]  ( .D(N120), .CLK(clk), .RSTB(n352), .Q(reg_b[28]) );
  DFFARX1 \reg_b_reg[18]  ( .D(N110), .CLK(clk), .RSTB(n347), .Q(reg_b[18]) );
  DFFARX1 \reg_b_reg[15]  ( .D(N107), .CLK(clk), .RSTB(n345), .Q(reg_b[15]) );
  DFFARX1 \reg_b_reg[9]  ( .D(N101), .CLK(clk), .RSTB(n342), .Q(reg_b[9]) );
  DFFARX1 \reg_b_reg[24]  ( .D(N116), .CLK(clk), .RSTB(n350), .Q(reg_b[24]) );
  DFFARX1 \reg_b_reg[26]  ( .D(N118), .CLK(clk), .RSTB(n351), .Q(reg_b[26]) );
  DFFARX1 \reg_b_reg[25]  ( .D(N117), .CLK(clk), .RSTB(n350), .Q(reg_b[25]) );
  DFFARX1 \reg_b_reg[27]  ( .D(N119), .CLK(clk), .RSTB(n351), .Q(reg_b[27]) );
  DFFARX1 \reg_b_reg[23]  ( .D(N115), .CLK(clk), .RSTB(n349), .Q(reg_b[23]) );
  DFFARX1 \reg_b_reg[13]  ( .D(N105), .CLK(clk), .RSTB(n344), .Q(reg_b[13]) );
  DFFARX1 \reg_b_reg[10]  ( .D(N102), .CLK(clk), .RSTB(n343), .Q(reg_b[10]), 
        .QN(n385) );
  DFFARX1 \reg_b_reg[30]  ( .D(N122), .CLK(clk), .RSTB(n353), .Q(reg_b[30]), 
        .QN(n554) );
  DFFARX1 \reg_b_reg[29]  ( .D(N121), .CLK(clk), .RSTB(n352), .Q(reg_b[29]), 
        .QN(n548) );
  DFFARX1 \reg_b_reg[19]  ( .D(N111), .CLK(clk), .RSTB(n347), .Q(reg_b[19]) );
  DFFARX1 \reg_b_reg[14]  ( .D(N106), .CLK(clk), .RSTB(n345), .Q(reg_b[14]) );
  DFFARX1 \reg_b_reg[20]  ( .D(N112), .CLK(clk), .RSTB(n348), .Q(reg_b[20]) );
  DFFARX1 \reg_b_reg[31]  ( .D(N123), .CLK(clk), .RSTB(n356), .Q(reg_b[31]), 
        .QN(n592) );
  DFFARX1 \reg_a_reg[19]  ( .D(N77), .CLK(clk), .RSTB(n347), .Q(reg_a[19]), 
        .QN(n392) );
  DFFARX1 \reg_a_reg[13]  ( .D(N71), .CLK(clk), .RSTB(n344), .Q(reg_a[13]), 
        .QN(n369) );
  DFFARX1 \reg_a_reg[22]  ( .D(N80), .CLK(clk), .RSTB(n349), .Q(reg_a[22]) );
  DFFARX1 \reg_a_reg[20]  ( .D(N78), .CLK(clk), .RSTB(n348), .Q(reg_a[20]), 
        .QN(n400) );
  DFFARX1 \reg_a_reg[9]  ( .D(N67), .CLK(clk), .RSTB(n342), .Q(reg_a[9]), .QN(
        n388) );
  DFFARX1 \reg_a_reg[31]  ( .D(N89), .CLK(clk), .RSTB(n357), .Q(reg_a[31]), 
        .QN(n430) );
  DFFARX1 \reg_a_reg[12]  ( .D(N70), .CLK(clk), .RSTB(n344), .Q(n113), .QN(
        n156) );
  DFFARX1 \reg_a_reg[25]  ( .D(N83), .CLK(clk), .RSTB(n350), .Q(reg_a[25]), 
        .QN(n417) );
  DFFARX1 \reg_a_reg[26]  ( .D(N84), .CLK(clk), .RSTB(n351), .Q(reg_a[26]), 
        .QN(n419) );
  DFFARX1 \reg_a_reg[27]  ( .D(N85), .CLK(clk), .RSTB(n351), .Q(reg_a[27]), 
        .QN(n424) );
  DFFARX1 \reg_a_reg[18]  ( .D(N76), .CLK(clk), .RSTB(n347), .Q(reg_a[18]), 
        .QN(n391) );
  DFFARX1 \reg_a_reg[23]  ( .D(N81), .CLK(clk), .RSTB(n349), .Q(reg_a[23]), 
        .QN(n411) );
  DFFARX1 \reg_a_reg[14]  ( .D(N72), .CLK(clk), .RSTB(n345), .Q(reg_a[14]), 
        .QN(n370) );
  DFFARX1 \reg_a_reg[28]  ( .D(N86), .CLK(clk), .RSTB(n352), .Q(reg_a[28]), 
        .QN(n427) );
  DFFARX1 \reg_a_reg[24]  ( .D(N82), .CLK(clk), .RSTB(n350), .Q(reg_a[24]), 
        .QN(n414) );
  DFFARX1 \reg_a_reg[6]  ( .D(N64), .CLK(clk), .RSTB(n355), .Q(reg_a[6]), .QN(
        n116) );
  DFFARX1 \reg_b_reg[12]  ( .D(N104), .CLK(clk), .RSTB(n344), .Q(reg_b[12]), 
        .QN(n213) );
  DFFARX1 \reg_b_reg[1]  ( .D(N93), .CLK(clk), .RSTB(n357), .Q(reg_b[1]), .QN(
        n241) );
  DFFARX1 \reg_a_reg[11]  ( .D(N69), .CLK(clk), .RSTB(n343), .Q(reg_a[11]), 
        .QN(n224) );
  DFFARX1 \reg_b_reg[4]  ( .D(N96), .CLK(clk), .RSTB(n354), .Q(reg_b[4]), .QN(
        n221) );
  DFFARX1 \reg_b_reg[11]  ( .D(N103), .CLK(clk), .RSTB(n343), .QN(n233) );
  DFFARX1 \reg_a_reg[4]  ( .D(N62), .CLK(clk), .RSTB(n354), .Q(reg_a[4]), .QN(
        n211) );
  DFFARX1 \reg_a_reg[15]  ( .D(N73), .CLK(clk), .RSTB(n345), .Q(reg_a[15]), 
        .QN(n145) );
  DFFARX1 \reg_a_reg[17]  ( .D(N75), .CLK(clk), .RSTB(n346), .Q(reg_a[17]), 
        .QN(n201) );
  DFFARX2 \reg_a_reg[8]  ( .D(N66), .CLK(clk), .RSTB(n342), .Q(reg_a[8]) );
  INVX4 U166 ( .IN(n480), .QN(n456) );
  XOR3X2 U167 ( .IN1(reg_b[26]), .IN2(reg_a[26]), .IN3(n538), .Q(n540) );
  NAND2X4 U168 ( .IN1(n413), .IN2(n135), .QN(n139) );
  OR2X4 U169 ( .IN1(n186), .IN2(n439), .Q(n596) );
  INVX2 U170 ( .IN(n187), .QN(n111) );
  XOR3X2 U171 ( .IN1(n201), .IN2(reg_b[17]), .IN3(n202), .Q(n492) );
  NAND2X4 U172 ( .IN1(n212), .IN2(reg_a[8]), .QN(n444) );
  INVX4 U173 ( .IN(reg_a[4]), .QN(n102) );
  INVX8 U174 ( .IN(n102), .QN(n103) );
  NOR2X4 U175 ( .IN1(n226), .IN2(n374), .QN(n376) );
  NAND2X2 U176 ( .IN1(n562), .IN2(n567), .QN(n374) );
  XOR3X2 U177 ( .IN1(reg_b[27]), .IN2(reg_a[27]), .IN3(n541), .Q(n543) );
  INVX4 U178 ( .IN(n541), .QN(n421) );
  NAND2X4 U179 ( .IN1(n138), .IN2(n459), .QN(n468) );
  NAND2X1 U180 ( .IN1(n224), .IN2(n258), .QN(n459) );
  INVX4 U181 ( .IN(reg_b[12]), .QN(n104) );
  INVX8 U182 ( .IN(n104), .QN(n105) );
  OR2X2 U183 ( .IN1(n382), .IN2(n229), .Q(n442) );
  INVX2 U184 ( .IN(n436), .QN(n382) );
  NAND2X2 U185 ( .IN1(n256), .IN2(n257), .QN(n454) );
  NAND2X1 U186 ( .IN1(n239), .IN2(reg_b[10]), .QN(n256) );
  INVX4 U187 ( .IN(n180), .QN(n181) );
  INVX4 U188 ( .IN(n188), .QN(n180) );
  XOR3X2 U189 ( .IN1(n103), .IN2(reg_b[4]), .IN3(n209), .Q(n574) );
  NAND2X2 U190 ( .IN1(n221), .IN2(n103), .QN(n576) );
  INVX8 U191 ( .IN(n123), .QN(n182) );
  OR2X4 U192 ( .IN1(n284), .IN2(n187), .Q(n123) );
  NAND2X2 U193 ( .IN1(n136), .IN2(n481), .QN(n195) );
  NAND2X0 U194 ( .IN1(reg_b[20]), .IN2(n400), .QN(n172) );
  INVX2 U195 ( .IN(n576), .QN(n378) );
  OAI21X1 U196 ( .IN1(reg_a[5]), .IN2(n215), .IN3(n575), .QN(n582) );
  INVX0 U197 ( .IN(n467), .QN(n372) );
  NAND2X0 U198 ( .IN1(reg_b[24]), .IN2(n414), .QN(n412) );
  OR2X1 U199 ( .IN1(reg_b[19]), .IN2(n392), .Q(n510) );
  INVX0 U200 ( .IN(n495), .QN(n394) );
  NOR2X0 U201 ( .IN1(reg_a[31]), .IN2(n592), .QN(n432) );
  NBUFFX2 U202 ( .IN(n119), .Q(n281) );
  NAND2X1 U203 ( .IN1(n207), .IN2(n581), .QN(n379) );
  NAND2X1 U204 ( .IN1(n582), .IN2(n581), .QN(n381) );
  NAND2X2 U205 ( .IN1(n393), .IN2(n397), .QN(n399) );
  NAND2X2 U206 ( .IN1(n192), .IN2(n450), .QN(n384) );
  OR4X1 U207 ( .IN1(reg_b[28]), .IN2(reg_b[29]), .IN3(reg_b[2]), .IN4(
        reg_b[30]), .Q(n60) );
  INVX2 U208 ( .IN(n529), .QN(n408) );
  OR2X1 U209 ( .IN1(reg_a[22]), .IN2(n225), .Q(n403) );
  NBUFFX2 U210 ( .IN(n442), .Q(n146) );
  NAND2X0 U211 ( .IN1(n220), .IN2(reg_a[21]), .QN(n524) );
  NAND2X0 U212 ( .IN1(n214), .IN2(reg_b[21]), .QN(n523) );
  INVX0 U213 ( .IN(n515), .QN(n517) );
  OAI21X1 U214 ( .IN1(reg_a[8]), .IN2(n212), .IN3(n435), .QN(n445) );
  OR2X1 U215 ( .IN1(n185), .IN2(n602), .Q(n562) );
  INVX0 U216 ( .IN(n241), .QN(n185) );
  NOR2X0 U217 ( .IN1(n613), .IN2(n284), .QN(n187) );
  NAND2X0 U218 ( .IN1(reg_b[28]), .IN2(n427), .QN(n425) );
  AND2X1 U219 ( .IN1(n207), .IN2(n580), .Q(n583) );
  NAND2X0 U220 ( .IN1(n153), .IN2(n154), .QN(n475) );
  NAND2X0 U221 ( .IN1(reg_b[13]), .IN2(n369), .QN(n154) );
  NAND2X1 U222 ( .IN1(n468), .IN2(n467), .QN(n153) );
  OR2X1 U223 ( .IN1(reg_b[13]), .IN2(n369), .Q(n474) );
  AND2X1 U224 ( .IN1(n473), .IN2(n480), .Q(n476) );
  NAND2X0 U225 ( .IN1(n210), .IN2(reg_a[17]), .QN(n495) );
  INVX0 U226 ( .IN(n493), .QN(n494) );
  INVX0 U227 ( .IN(n508), .QN(n509) );
  XOR3X1 U228 ( .IN1(reg_a[13]), .IN2(reg_b[13]), .IN3(n470), .Q(n471) );
  AND2X1 U229 ( .IN1(n466), .IN2(n480), .Q(n469) );
  INVX0 U230 ( .IN(n501), .QN(n502) );
  INVX0 U231 ( .IN(n435), .QN(n437) );
  INVX0 U232 ( .IN(n150), .QN(n491) );
  AND2X1 U233 ( .IN1(n136), .IN2(n480), .Q(n483) );
  INVX0 U234 ( .IN(n147), .QN(n148) );
  NBUFFX8 U235 ( .IN(n119), .Q(n284) );
  NOR2X0 U236 ( .IN1(reg_b[31]), .IN2(n430), .QN(n431) );
  INVX0 U237 ( .IN(n116), .QN(n236) );
  INVX2 U238 ( .IN(n434), .QN(n613) );
  INVX2 U239 ( .IN(n106), .QN(n107) );
  INVX2 U240 ( .IN(reg_a[7]), .QN(n106) );
  INVX0 U241 ( .IN(n173), .QN(n532) );
  INVX0 U242 ( .IN(n167), .QN(n544) );
  XOR3X1 U243 ( .IN1(reg_b[23]), .IN2(reg_a[23]), .IN3(n529), .Q(n531) );
  XOR3X1 U244 ( .IN1(reg_b[25]), .IN2(reg_a[25]), .IN3(n535), .Q(n537) );
  NOR2X0 U245 ( .IN1(n416), .IN2(n415), .QN(n535) );
  XOR3X1 U246 ( .IN1(n113), .IN2(n105), .IN3(n462), .Q(n464) );
  NAND2X0 U247 ( .IN1(n267), .IN2(n268), .QN(n593) );
  NAND2X0 U248 ( .IN1(b_in[18]), .IN2(n281), .QN(n170) );
  NAND2X0 U249 ( .IN1(n275), .IN2(reg_b[18]), .QN(n168) );
  XOR3X1 U250 ( .IN1(n237), .IN2(reg_b[2]), .IN3(n194), .Q(n565) );
  XOR3X1 U251 ( .IN1(reg_a[16]), .IN2(n262), .IN3(n193), .Q(n490) );
  XOR3X1 U252 ( .IN1(reg_b[10]), .IN2(reg_a[10]), .IN3(n453), .Q(n455) );
  NAND2X0 U253 ( .IN1(n606), .IN2(n605), .QN(N59) );
  NOR2X0 U254 ( .IN1(n600), .IN2(n599), .QN(n606) );
  INVX0 U255 ( .IN(n413), .QN(n416) );
  NAND2X4 U256 ( .IN1(n412), .IN2(n173), .QN(n413) );
  NAND2X4 U257 ( .IN1(n428), .IN2(n155), .QN(n222) );
  NAND2X2 U258 ( .IN1(n496), .IN2(n495), .QN(n259) );
  NAND2X2 U259 ( .IN1(n511), .IN2(n510), .QN(n171) );
  OR4X2 U260 ( .IN1(reg_b[17]), .IN2(reg_b[18]), .IN3(reg_b[19]), .IN4(
        reg_b[1]), .Q(n63) );
  NAND2X4 U261 ( .IN1(n377), .IN2(n566), .QN(n580) );
  AND2X2 U262 ( .IN1(n426), .IN2(n115), .Q(n557) );
  NAND2X4 U263 ( .IN1(n167), .IN2(n425), .QN(n426) );
  NAND2X4 U264 ( .IN1(n139), .IN2(n121), .QN(n538) );
  OR4X4 U265 ( .IN1(reg_b[13]), .IN2(reg_b[14]), .IN3(reg_b[15]), .IN4(n262), 
        .Q(n64) );
  NOR2X0 U266 ( .IN1(n262), .IN2(n216), .QN(n150) );
  AND2X2 U267 ( .IN1(n216), .IN2(n262), .Q(n124) );
  INVX4 U268 ( .IN(n261), .QN(n262) );
  NOR2X4 U269 ( .IN1(n380), .IN2(n175), .QN(n174) );
  INVX4 U270 ( .IN(n596), .QN(n108) );
  INVX4 U271 ( .IN(n596), .QN(n109) );
  INVX1 U272 ( .IN(n186), .QN(n110) );
  NAND2X0 U273 ( .IN1(n199), .IN2(n200), .QN(n6) );
  OR2X1 U274 ( .IN1(n236), .IN2(n230), .Q(n112) );
  AND2X1 U275 ( .IN1(n227), .IN2(n100), .Q(n114) );
  OR2X1 U276 ( .IN1(reg_b[28]), .IN2(n427), .Q(n115) );
  OR2X1 U277 ( .IN1(reg_b[23]), .IN2(n411), .Q(n117) );
  OR2X1 U278 ( .IN1(reg_b[27]), .IN2(n424), .Q(n118) );
  NAND2X2 U279 ( .IN1(n259), .IN2(n260), .QN(n504) );
  AND3X2 U280 ( .IN1(start), .IN2(n67), .IN3(n100), .Q(n119) );
  NOR2X0 U281 ( .IN1(n429), .IN2(n432), .QN(n120) );
  NAND2X0 U282 ( .IN1(n140), .IN2(n157), .QN(n121) );
  NOR2X0 U283 ( .IN1(n368), .IN2(n141), .QN(n122) );
  NBUFFX2 U284 ( .IN(n572), .Q(n143) );
  INVX2 U285 ( .IN(n519), .QN(n397) );
  NAND2X2 U286 ( .IN1(n171), .IN2(n172), .QN(n519) );
  AOI22X1 U287 ( .IN1(n239), .IN2(reg_b[9]), .IN3(n166), .IN4(reg_a[9]), .QN(
        n125) );
  AOI22X1 U288 ( .IN1(n239), .IN2(reg_b[13]), .IN3(n165), .IN4(reg_a[13]), 
        .QN(n126) );
  AOI22X1 U289 ( .IN1(n239), .IN2(reg_b[20]), .IN3(n166), .IN4(reg_a[20]), 
        .QN(n127) );
  AOI22X1 U290 ( .IN1(n239), .IN2(reg_b[8]), .IN3(n165), .IN4(reg_a[8]), .QN(
        n128) );
  AOI22X1 U291 ( .IN1(n239), .IN2(reg_b[19]), .IN3(n165), .IN4(reg_a[19]), 
        .QN(n129) );
  AOI22X1 U292 ( .IN1(n239), .IN2(reg_b[22]), .IN3(n165), .IN4(reg_a[22]), 
        .QN(n130) );
  AOI22X1 U293 ( .IN1(n239), .IN2(reg_b[6]), .IN3(n165), .IN4(n236), .QN(n131)
         );
  AOI22X1 U294 ( .IN1(n239), .IN2(reg_b[21]), .IN3(n165), .IN4(reg_a[21]), 
        .QN(n132) );
  AOI22X1 U295 ( .IN1(n239), .IN2(reg_b[17]), .IN3(n166), .IN4(reg_a[17]), 
        .QN(n133) );
  AOI22X1 U296 ( .IN1(n239), .IN2(reg_b[5]), .IN3(n166), .IN4(n148), .QN(n134)
         );
  NOR2X0 U297 ( .IN1(n415), .IN2(n418), .QN(n135) );
  INVX0 U298 ( .IN(n178), .QN(n179) );
  NOR2X0 U299 ( .IN1(n373), .IN2(n472), .QN(n136) );
  AND2X1 U300 ( .IN1(n122), .IN2(n115), .Q(n137) );
  OR2X2 U301 ( .IN1(n205), .IN2(n487), .Q(n516) );
  NAND2X2 U302 ( .IN1(n156), .IN2(n105), .QN(n138) );
  NAND2X4 U303 ( .IN1(n482), .IN2(n481), .QN(n217) );
  NAND2X0 U304 ( .IN1(n222), .IN2(n223), .QN(n588) );
  OR4X4 U305 ( .IN1(n176), .IN2(reg_b[10]), .IN3(n258), .IN4(n105), .Q(n65) );
  INVX0 U306 ( .IN(n418), .QN(n140) );
  INVX0 U307 ( .IN(n555), .QN(n141) );
  NAND2X4 U308 ( .IN1(n137), .IN2(n426), .QN(n428) );
  NAND2X4 U309 ( .IN1(n222), .IN2(n142), .QN(n434) );
  AND2X1 U310 ( .IN1(n223), .IN2(n114), .Q(n142) );
  NAND2X4 U311 ( .IN1(n144), .IN2(reg_b[7]), .QN(n435) );
  AO21X1 U312 ( .IN1(n201), .IN2(reg_b[17]), .IN3(n124), .Q(n496) );
  INVX4 U313 ( .IN(n580), .QN(n572) );
  OR2X2 U314 ( .IN1(n372), .IN2(n465), .Q(n472) );
  OR2X2 U315 ( .IN1(n231), .IN2(n371), .Q(n465) );
  NOR2X4 U316 ( .IN1(reg_b[10]), .IN2(n196), .QN(n231) );
  INVX0 U317 ( .IN(n449), .QN(n149) );
  NOR2X4 U318 ( .IN1(n378), .IN2(n228), .QN(n207) );
  NOR2X4 U319 ( .IN1(n442), .IN2(n383), .QN(n192) );
  NAND2X4 U320 ( .IN1(n397), .IN2(n515), .QN(n398) );
  OR2X2 U321 ( .IN1(n237), .IN2(n219), .Q(n566) );
  NAND2X0 U322 ( .IN1(n611), .IN2(n471), .QN(n151) );
  NAND2X0 U323 ( .IN1(a_in[13]), .IN2(n191), .QN(n152) );
  NAND3X0 U324 ( .IN1(n151), .IN2(n152), .IN3(n126), .QN(N71) );
  OR2X2 U325 ( .IN1(n396), .IN2(n508), .Q(n515) );
  INVX16 U326 ( .IN(n601), .QN(n166) );
  INVX8 U327 ( .IN(n163), .QN(n601) );
  NOR2X4 U328 ( .IN1(n376), .IN2(n375), .QN(n377) );
  NAND2X2 U329 ( .IN1(n213), .IN2(n113), .QN(n467) );
  AND2X1 U330 ( .IN1(n553), .IN2(n120), .Q(n155) );
  AND2X2 U331 ( .IN1(n230), .IN2(reg_a[6]), .Q(n229) );
  NAND2X1 U332 ( .IN1(n239), .IN2(reg_b[31]), .QN(n267) );
  NOR2X4 U333 ( .IN1(n387), .IN2(n386), .QN(n390) );
  NOR2X4 U334 ( .IN1(n174), .IN2(n384), .QN(n387) );
  NAND2X2 U335 ( .IN1(n240), .IN2(n107), .QN(n436) );
  AND2X1 U336 ( .IN1(reg_b[25]), .IN2(n417), .Q(n157) );
  NOR2X4 U337 ( .IN1(n538), .IN2(n159), .QN(n158) );
  AND2X1 U338 ( .IN1(reg_b[26]), .IN2(n419), .Q(n159) );
  AND2X4 U339 ( .IN1(n192), .IN2(n449), .Q(n452) );
  INVX8 U340 ( .IN(n597), .QN(n160) );
  INVX8 U341 ( .IN(n597), .QN(n611) );
  NAND2X4 U342 ( .IN1(n445), .IN2(n444), .QN(n161) );
  NAND2X4 U343 ( .IN1(reg_b[9]), .IN2(n388), .QN(n162) );
  NAND2X4 U344 ( .IN1(n161), .IN2(n162), .QN(n451) );
  NAND2X4 U345 ( .IN1(n451), .IN2(n450), .QN(n389) );
  NOR2X4 U346 ( .IN1(n440), .IN2(n110), .QN(n163) );
  INVX8 U347 ( .IN(n271), .QN(n238) );
  NOR2X4 U348 ( .IN1(n203), .IN2(n440), .QN(n271) );
  INVX2 U349 ( .IN(n221), .QN(n164) );
  NOR2X4 U350 ( .IN1(n613), .IN2(n284), .QN(n186) );
  INVX8 U351 ( .IN(n601), .QN(n165) );
  NAND2X4 U352 ( .IN1(n423), .IN2(n118), .QN(n167) );
  NAND2X0 U353 ( .IN1(n182), .IN2(reg_a[18]), .QN(n169) );
  NAND3X0 U354 ( .IN1(n168), .IN2(n169), .IN3(n170), .QN(N110) );
  NAND2X4 U355 ( .IN1(n410), .IN2(n117), .QN(n173) );
  IBUFFX16 U356 ( .IN(n174), .QN(n449) );
  NAND2X2 U357 ( .IN1(n381), .IN2(n112), .QN(n175) );
  NOR2X4 U358 ( .IN1(n572), .IN2(n379), .QN(n380) );
  NOR2X0 U359 ( .IN1(n613), .IN2(n284), .QN(n177) );
  INVX2 U360 ( .IN(n234), .QN(n183) );
  NOR2X0 U361 ( .IN1(n613), .IN2(n284), .QN(n203) );
  DELLN3X2 U362 ( .IN(reg_a[1]), .Q(n184) );
  INVX32 U363 ( .IN(n238), .QN(n239) );
  NOR2X2 U364 ( .IN1(n284), .IN2(n186), .QN(n188) );
  NBUFFX2 U365 ( .IN(n613), .Q(n190) );
  NOR2X0 U366 ( .IN1(n368), .IN2(n547), .QN(n429) );
  NOR2X0 U367 ( .IN1(reg_b[3]), .IN2(n235), .QN(n228) );
  NAND2X1 U368 ( .IN1(n211), .IN2(n164), .QN(n575) );
  INVX4 U369 ( .IN(n596), .QN(n191) );
  INVX4 U370 ( .IN(n596), .QN(n609) );
  OR2X2 U371 ( .IN1(n150), .IN2(n232), .Q(n493) );
  INVX2 U372 ( .IN(n460), .QN(n371) );
  OR2X2 U373 ( .IN1(n395), .IN2(n501), .Q(n508) );
  NAND2X4 U374 ( .IN1(n524), .IN2(n518), .QN(n401) );
  NOR2X0 U375 ( .IN1(n232), .IN2(n488), .QN(n193) );
  NOR2X0 U376 ( .IN1(n226), .IN2(n563), .QN(n194) );
  AND2X1 U377 ( .IN1(n225), .IN2(reg_a[22]), .Q(n406) );
  NOR2X0 U378 ( .IN1(reg_a[10]), .IN2(n385), .QN(n386) );
  OR2X1 U379 ( .IN1(reg_b[18]), .IN2(n391), .Q(n503) );
  NAND2X0 U380 ( .IN1(reg_b[15]), .IN2(n145), .QN(n218) );
  OR2X1 U381 ( .IN1(reg_b[30]), .IN2(n197), .Q(n589) );
  OR2X1 U382 ( .IN1(reg_b[29]), .IN2(n198), .Q(n555) );
  NAND2X2 U383 ( .IN1(reg_b[23]), .IN2(n411), .QN(n409) );
  NAND2X1 U384 ( .IN1(reg_b[27]), .IN2(n424), .QN(n422) );
  NAND2X0 U385 ( .IN1(n163), .IN2(reg_a[10]), .QN(n257) );
  XOR3X1 U386 ( .IN1(n184), .IN2(n607), .IN3(reg_b[1]), .Q(n598) );
  NOR4X0 U387 ( .IN1(n64), .IN2(n65), .IN3(n62), .IN4(n63), .QN(n199) );
  NOR4X0 U388 ( .IN1(n60), .IN2(n61), .IN3(n58), .IN4(n59), .QN(n200) );
  NOR2X0 U389 ( .IN1(n100), .IN2(n227), .QN(done) );
  OAI21X1 U390 ( .IN1(n124), .IN2(n193), .IN3(n491), .QN(n202) );
  NAND2X2 U391 ( .IN1(n270), .IN2(n183), .QN(n607) );
  NOR2X4 U392 ( .IN1(n456), .IN2(n195), .QN(n205) );
  INVX0 U393 ( .IN(n324), .QN(n306) );
  INVX0 U394 ( .IN(n324), .QN(n305) );
  INVX0 U395 ( .IN(n326), .QN(n302) );
  INVX0 U396 ( .IN(n320), .QN(n314) );
  INVX0 U397 ( .IN(n320), .QN(n313) );
  INVX0 U398 ( .IN(n321), .QN(n312) );
  INVX0 U399 ( .IN(n321), .QN(n311) );
  INVX0 U400 ( .IN(n322), .QN(n310) );
  INVX0 U401 ( .IN(n322), .QN(n309) );
  INVX0 U402 ( .IN(n323), .QN(n308) );
  INVX0 U403 ( .IN(n323), .QN(n307) );
  INVX0 U404 ( .IN(n325), .QN(n304) );
  INVX0 U405 ( .IN(n325), .QN(n303) );
  INVX0 U406 ( .IN(n285), .QN(n320) );
  INVX0 U407 ( .IN(n285), .QN(n321) );
  INVX0 U408 ( .IN(n286), .QN(n322) );
  INVX0 U409 ( .IN(n286), .QN(n323) );
  INVX0 U410 ( .IN(n287), .QN(n324) );
  INVX0 U411 ( .IN(n287), .QN(n325) );
  INVX0 U412 ( .IN(n288), .QN(n326) );
  INVX0 U413 ( .IN(n295), .QN(n341) );
  INVX0 U414 ( .IN(n295), .QN(n340) );
  INVX0 U415 ( .IN(n294), .QN(n339) );
  INVX0 U416 ( .IN(n294), .QN(n338) );
  INVX0 U417 ( .IN(n293), .QN(n337) );
  INVX0 U418 ( .IN(n293), .QN(n336) );
  INVX0 U419 ( .IN(n292), .QN(n335) );
  INVX0 U420 ( .IN(n291), .QN(n333) );
  INVX0 U421 ( .IN(n291), .QN(n332) );
  INVX0 U422 ( .IN(n290), .QN(n331) );
  INVX0 U423 ( .IN(n289), .QN(n328) );
  INVX0 U424 ( .IN(n288), .QN(n327) );
  INVX0 U425 ( .IN(n292), .QN(n334) );
  INVX0 U426 ( .IN(n290), .QN(n330) );
  INVX0 U427 ( .IN(n289), .QN(n329) );
  INVX0 U428 ( .IN(n299), .QN(n317) );
  INVX0 U429 ( .IN(n319), .QN(n316) );
  INVX0 U430 ( .IN(n319), .QN(n315) );
  INVX0 U431 ( .IN(n301), .QN(n318) );
  INVX0 U432 ( .IN(n301), .QN(n285) );
  INVX0 U433 ( .IN(n301), .QN(n286) );
  INVX0 U434 ( .IN(n300), .QN(n287) );
  INVX0 U435 ( .IN(n300), .QN(n288) );
  INVX0 U436 ( .IN(n296), .QN(n295) );
  INVX0 U437 ( .IN(n295), .QN(n319) );
  INVX0 U438 ( .IN(n297), .QN(n294) );
  INVX0 U439 ( .IN(n297), .QN(n293) );
  INVX0 U440 ( .IN(n298), .QN(n291) );
  INVX0 U441 ( .IN(n299), .QN(n290) );
  INVX0 U442 ( .IN(n299), .QN(n289) );
  INVX0 U443 ( .IN(n298), .QN(n292) );
  AND2X1 U444 ( .IN1(n114), .IN2(n318), .Q(n433) );
  OR3X1 U445 ( .IN1(n190), .IN2(n612), .IN3(n276), .Q(gcd_ns[0]) );
  AND2X1 U446 ( .IN1(n114), .IN2(n318), .Q(n612) );
  AND2X1 U447 ( .IN1(n494), .IN2(n516), .Q(n497) );
  NOR2X0 U448 ( .IN1(n456), .IN2(n231), .QN(n204) );
  INVX0 U449 ( .IN(n6), .QN(n301) );
  INVX0 U450 ( .IN(n6), .QN(n300) );
  INVX0 U451 ( .IN(n6), .QN(n297) );
  INVX0 U452 ( .IN(n6), .QN(n299) );
  INVX0 U453 ( .IN(n6), .QN(n296) );
  INVX0 U454 ( .IN(n6), .QN(n298) );
  INVX0 U455 ( .IN(n510), .QN(n396) );
  NOR2X0 U456 ( .IN1(n604), .IN2(n603), .QN(n605) );
  NOR2X0 U457 ( .IN1(n596), .IN2(n595), .QN(n600) );
  INVX0 U458 ( .IN(n444), .QN(n383) );
  INVX0 U459 ( .IN(n503), .QN(n395) );
  OR2X2 U460 ( .IN1(n394), .IN2(n493), .Q(n501) );
  INVX0 U461 ( .IN(n474), .QN(n373) );
  INVX0 U462 ( .IN(n465), .QN(n466) );
  INVX0 U463 ( .IN(n472), .QN(n473) );
  INVX0 U464 ( .IN(n589), .QN(n368) );
  OA21X1 U465 ( .IN1(n557), .IN2(n556), .IN3(n555), .Q(n206) );
  NBUFFX2 U466 ( .IN(n119), .Q(n279) );
  NBUFFX2 U467 ( .IN(n119), .Q(n276) );
  NBUFFX2 U468 ( .IN(n119), .Q(n282) );
  NBUFFX2 U469 ( .IN(n119), .Q(n280) );
  NBUFFX2 U470 ( .IN(n119), .Q(n278) );
  NBUFFX2 U471 ( .IN(n119), .Q(n283) );
  NBUFFX2 U472 ( .IN(n119), .Q(n277) );
  INVX0 U473 ( .IN(n459), .QN(n461) );
  OR2X1 U474 ( .IN1(n368), .IN2(n590), .Q(n559) );
  INVX0 U475 ( .IN(n521), .QN(n525) );
  AND2X1 U476 ( .IN1(n517), .IN2(n516), .Q(n520) );
  NOR2X0 U477 ( .IN1(n149), .IN2(n229), .QN(n208) );
  NOR2X0 U478 ( .IN1(n143), .IN2(n228), .QN(n209) );
  INVX0 U479 ( .IN(n547), .QN(n556) );
  INVX0 U480 ( .IN(n553), .QN(n590) );
  INVX0 U481 ( .IN(n562), .QN(n563) );
  INVX0 U482 ( .IN(n516), .QN(n488) );
  OR2X1 U483 ( .IN1(n141), .IN2(n556), .Q(n550) );
  INVX0 U484 ( .IN(n566), .QN(n568) );
  NBUFFX2 U485 ( .IN(n359), .Q(n357) );
  NBUFFX2 U486 ( .IN(n364), .Q(n347) );
  NBUFFX2 U487 ( .IN(n361), .Q(n353) );
  NBUFFX2 U488 ( .IN(n360), .Q(n356) );
  NBUFFX2 U489 ( .IN(n366), .Q(n343) );
  NBUFFX2 U490 ( .IN(n366), .Q(n344) );
  NBUFFX2 U491 ( .IN(n365), .Q(n346) );
  NBUFFX2 U492 ( .IN(n364), .Q(n348) );
  NBUFFX2 U493 ( .IN(n362), .Q(n352) );
  NBUFFX2 U494 ( .IN(n360), .Q(n355) );
  NBUFFX2 U495 ( .IN(n365), .Q(n345) );
  NBUFFX2 U496 ( .IN(n363), .Q(n349) );
  NBUFFX2 U497 ( .IN(n363), .Q(n350) );
  NBUFFX2 U498 ( .IN(n362), .Q(n351) );
  NBUFFX2 U499 ( .IN(n361), .Q(n354) );
  NBUFFX2 U500 ( .IN(n359), .Q(n358) );
  NAND2X0 U501 ( .IN1(n163), .IN2(reg_a[31]), .QN(n268) );
  OR2X1 U502 ( .IN1(reg_b[14]), .IN2(n370), .Q(n481) );
  NAND2X0 U503 ( .IN1(a_in[21]), .IN2(n191), .QN(n253) );
  OR2X1 U504 ( .IN1(n258), .IN2(n224), .Q(n460) );
  AO222X1 U505 ( .IN1(n275), .IN2(reg_b[13]), .IN3(n181), .IN4(reg_a[13]), 
        .IN5(b_in[13]), .IN6(n282), .Q(N105) );
  AO222X1 U506 ( .IN1(n275), .IN2(reg_b[14]), .IN3(n181), .IN4(reg_a[14]), 
        .IN5(b_in[14]), .IN6(n282), .Q(N106) );
  AO222X1 U507 ( .IN1(n272), .IN2(reg_b[19]), .IN3(n181), .IN4(reg_a[19]), 
        .IN5(b_in[19]), .IN6(n281), .Q(N111) );
  AO222X1 U508 ( .IN1(n274), .IN2(reg_b[23]), .IN3(n181), .IN4(reg_a[23]), 
        .IN5(b_in[23]), .IN6(n280), .Q(N115) );
  AO222X1 U509 ( .IN1(n275), .IN2(reg_b[25]), .IN3(n181), .IN4(reg_a[25]), 
        .IN5(b_in[25]), .IN6(n279), .Q(N117) );
  AO222X1 U510 ( .IN1(n272), .IN2(reg_b[26]), .IN3(n181), .IN4(reg_a[26]), 
        .IN5(b_in[26]), .IN6(n279), .Q(N118) );
  AO222X1 U511 ( .IN1(n273), .IN2(reg_b[27]), .IN3(n181), .IN4(reg_a[27]), 
        .IN5(b_in[27]), .IN6(n279), .Q(N119) );
  AO222X1 U512 ( .IN1(n273), .IN2(reg_b[8]), .IN3(n181), .IN4(reg_a[8]), .IN5(
        b_in[8]), .IN6(n284), .Q(N100) );
  AO222X1 U513 ( .IN1(n272), .IN2(n105), .IN3(n181), .IN4(n113), .IN5(b_in[12]), .IN6(n283), .Q(N104) );
  AO222X1 U514 ( .IN1(n272), .IN2(reg_b[17]), .IN3(n188), .IN4(reg_a[17]), 
        .IN5(b_in[17]), .IN6(n281), .Q(N109) );
  AO222X1 U515 ( .IN1(n272), .IN2(reg_b[5]), .IN3(n188), .IN4(n148), .IN5(
        b_in[5]), .IN6(n277), .Q(N97) );
  AO222X1 U516 ( .IN1(n272), .IN2(reg_b[21]), .IN3(n188), .IN4(reg_a[21]), 
        .IN5(b_in[21]), .IN6(n280), .Q(N113) );
  AO222X1 U517 ( .IN1(n275), .IN2(reg_b[20]), .IN3(n181), .IN4(reg_a[20]), 
        .IN5(b_in[20]), .IN6(n281), .Q(N112) );
  AO222X1 U518 ( .IN1(n274), .IN2(reg_b[29]), .IN3(n188), .IN4(reg_a[29]), 
        .IN5(b_in[29]), .IN6(n278), .Q(N121) );
  AO222X1 U519 ( .IN1(n274), .IN2(reg_b[30]), .IN3(n188), .IN4(reg_a[30]), 
        .IN5(b_in[30]), .IN6(n278), .Q(N122) );
  OR4X1 U520 ( .IN1(reg_b[20]), .IN2(reg_b[21]), .IN3(reg_b[22]), .IN4(
        reg_b[23]), .Q(n62) );
  OR4X1 U521 ( .IN1(reg_b[24]), .IN2(reg_b[25]), .IN3(reg_b[26]), .IN4(
        reg_b[27]), .Q(n61) );
  OR2X1 U522 ( .IN1(reg_a[29]), .IN2(n548), .Q(n547) );
  OR2X1 U523 ( .IN1(reg_a[30]), .IN2(n554), .Q(n553) );
  AND2X1 U524 ( .IN1(reg_b[1]), .IN2(n239), .Q(n603) );
  AO22X1 U525 ( .IN1(reg_a[8]), .IN2(n339), .IN3(result[8]), .IN4(n317), .Q(
        n68) );
  AO22X1 U526 ( .IN1(reg_a[9]), .IN2(n341), .IN3(result[9]), .IN4(n317), .Q(
        n69) );
  AO22X1 U527 ( .IN1(reg_a[10]), .IN2(n341), .IN3(result[10]), .IN4(n316), .Q(
        n70) );
  AO22X1 U528 ( .IN1(reg_a[11]), .IN2(n340), .IN3(result[11]), .IN4(n316), .Q(
        n71) );
  AO22X1 U529 ( .IN1(n113), .IN2(n340), .IN3(result[12]), .IN4(n315), .Q(n72)
         );
  AO22X1 U530 ( .IN1(reg_a[13]), .IN2(n339), .IN3(result[13]), .IN4(n315), .Q(
        n73) );
  AO22X1 U531 ( .IN1(reg_a[14]), .IN2(n339), .IN3(result[14]), .IN4(n314), .Q(
        n74) );
  AO22X1 U532 ( .IN1(reg_a[15]), .IN2(n338), .IN3(result[15]), .IN4(n314), .Q(
        n75) );
  AO22X1 U533 ( .IN1(reg_a[16]), .IN2(n338), .IN3(result[16]), .IN4(n313), .Q(
        n76) );
  AO22X1 U534 ( .IN1(reg_a[17]), .IN2(n337), .IN3(result[17]), .IN4(n313), .Q(
        n77) );
  AO22X1 U535 ( .IN1(reg_a[18]), .IN2(n337), .IN3(result[18]), .IN4(n312), .Q(
        n78) );
  AO22X1 U536 ( .IN1(reg_a[19]), .IN2(n336), .IN3(result[19]), .IN4(n312), .Q(
        n79) );
  AO22X1 U537 ( .IN1(reg_a[20]), .IN2(n336), .IN3(result[20]), .IN4(n311), .Q(
        n80) );
  AO22X1 U538 ( .IN1(reg_a[21]), .IN2(n335), .IN3(result[21]), .IN4(n311), .Q(
        n81) );
  AO22X1 U539 ( .IN1(reg_a[22]), .IN2(n335), .IN3(result[22]), .IN4(n310), .Q(
        n82) );
  AO22X1 U540 ( .IN1(reg_a[23]), .IN2(n334), .IN3(result[23]), .IN4(n310), .Q(
        n83) );
  AO22X1 U541 ( .IN1(reg_a[24]), .IN2(n333), .IN3(result[24]), .IN4(n309), .Q(
        n84) );
  AO22X1 U542 ( .IN1(reg_a[25]), .IN2(n333), .IN3(result[25]), .IN4(n309), .Q(
        n85) );
  AO22X1 U543 ( .IN1(reg_a[26]), .IN2(n332), .IN3(result[26]), .IN4(n308), .Q(
        n86) );
  AO22X1 U544 ( .IN1(reg_a[27]), .IN2(n332), .IN3(result[27]), .IN4(n308), .Q(
        n87) );
  AO22X1 U545 ( .IN1(reg_a[28]), .IN2(n331), .IN3(result[28]), .IN4(n307), .Q(
        n88) );
  AO22X1 U546 ( .IN1(reg_a[29]), .IN2(n331), .IN3(result[29]), .IN4(n307), .Q(
        n89) );
  AO22X1 U547 ( .IN1(reg_a[30]), .IN2(n330), .IN3(result[30]), .IN4(n306), .Q(
        n90) );
  AO22X1 U548 ( .IN1(reg_a[3]), .IN2(n329), .IN3(result[3]), .IN4(n305), .Q(
        n92) );
  AO22X1 U549 ( .IN1(n148), .IN2(n328), .IN3(result[5]), .IN4(n304), .Q(n94)
         );
  AO22X1 U550 ( .IN1(n236), .IN2(n328), .IN3(result[6]), .IN4(n304), .Q(n95)
         );
  AO22X1 U551 ( .IN1(n107), .IN2(n327), .IN3(result[7]), .IN4(n303), .Q(n96)
         );
  AO22X1 U552 ( .IN1(reg_a[31]), .IN2(n327), .IN3(result[31]), .IN4(n303), .Q(
        n97) );
  AO22X1 U553 ( .IN1(reg_a[0]), .IN2(n334), .IN3(result[0]), .IN4(n302), .Q(
        n99) );
  AND2X1 U554 ( .IN1(n184), .IN2(n166), .Q(n604) );
  XOR3X1 U555 ( .IN1(n107), .IN2(reg_b[7]), .IN3(n208), .Q(n587) );
  MUX21X1 U556 ( .IN1(n559), .IN2(n558), .S(n206), .Q(n561) );
  XOR2X1 U557 ( .IN1(n554), .IN2(reg_a[30]), .Q(n558) );
  XOR2X1 U558 ( .IN1(n548), .IN2(reg_a[29]), .Q(n549) );
  OA21X1 U559 ( .IN1(n461), .IN2(n204), .IN3(n460), .Q(n462) );
  OAI21X1 U560 ( .IN1(n176), .IN2(n270), .IN3(n607), .QN(n610) );
  AND3X1 U561 ( .IN1(reg_a[31]), .IN2(n592), .IN3(n591), .Q(n594) );
  OAI21X1 U562 ( .IN1(n590), .IN2(n206), .IN3(n589), .QN(n591) );
  OA21X1 U563 ( .IN1(n452), .IN2(n451), .IN3(n450), .Q(n453) );
  NAND2X2 U564 ( .IN1(n215), .IN2(n148), .QN(n581) );
  NOR2X0 U565 ( .IN1(n598), .IN2(n597), .QN(n599) );
  XOR3X1 U566 ( .IN1(reg_a[18]), .IN2(reg_b[18]), .IN3(n498), .Q(n500) );
  OA21X1 U567 ( .IN1(n497), .IN2(n496), .IN3(n495), .Q(n498) );
  XOR3X1 U568 ( .IN1(reg_a[14]), .IN2(reg_b[14]), .IN3(n477), .Q(n479) );
  XOR3X1 U569 ( .IN1(reg_b[28]), .IN2(reg_a[28]), .IN3(n544), .Q(n546) );
  XOR3X1 U570 ( .IN1(reg_b[24]), .IN2(reg_a[24]), .IN3(n532), .Q(n534) );
  XOR3X1 U571 ( .IN1(reg_a[11]), .IN2(n258), .IN3(n204), .Q(n458) );
  XOR3X1 U572 ( .IN1(reg_a[15]), .IN2(reg_b[15]), .IN3(n484), .Q(n486) );
  XOR3X1 U573 ( .IN1(n179), .IN2(reg_a[3]), .IN3(n569), .Q(n571) );
  OA21X1 U574 ( .IN1(n568), .IN2(n194), .IN3(n567), .Q(n569) );
  INVX4 U575 ( .IN(n233), .QN(n258) );
  NOR2X1 U576 ( .IN1(reg_a[3]), .IN2(n178), .QN(n375) );
  NAND2X4 U577 ( .IN1(n217), .IN2(n218), .QN(n487) );
  XOR3X1 U578 ( .IN1(reg_a[9]), .IN2(reg_b[9]), .IN3(n447), .Q(n448) );
  OA21X1 U579 ( .IN1(n446), .IN2(n445), .IN3(n444), .Q(n447) );
  AND2X1 U580 ( .IN1(n443), .IN2(n449), .Q(n446) );
  INVX0 U581 ( .IN(n146), .QN(n443) );
  XOR3X1 U582 ( .IN1(reg_a[19]), .IN2(reg_b[19]), .IN3(n506), .Q(n507) );
  AND2X1 U583 ( .IN1(n502), .IN2(n516), .Q(n505) );
  XOR3X1 U584 ( .IN1(reg_a[8]), .IN2(reg_b[8]), .IN3(n438), .Q(n441) );
  OA21X1 U585 ( .IN1(n437), .IN2(n208), .IN3(n436), .Q(n438) );
  XOR3X1 U586 ( .IN1(reg_a[21]), .IN2(reg_b[21]), .IN3(n525), .Q(n522) );
  XOR3X1 U587 ( .IN1(n148), .IN2(reg_b[5]), .IN3(n578), .Q(n579) );
  INVX0 U588 ( .IN(n575), .QN(n577) );
  NAND2X1 U589 ( .IN1(n219), .IN2(n237), .QN(n567) );
  XOR3X1 U590 ( .IN1(reg_b[20]), .IN2(reg_a[20]), .IN3(n513), .Q(n514) );
  AND2X1 U591 ( .IN1(n509), .IN2(n516), .Q(n512) );
  XOR3X1 U592 ( .IN1(reg_b[22]), .IN2(reg_a[22]), .IN3(n527), .Q(n528) );
  OA21X1 U593 ( .IN1(n526), .IN2(n525), .IN3(n524), .Q(n527) );
  INVX0 U594 ( .IN(n523), .QN(n526) );
  XOR3X1 U595 ( .IN1(reg_b[6]), .IN2(n236), .IN3(n584), .Q(n585) );
  OA21X1 U596 ( .IN1(n583), .IN2(n582), .IN3(n581), .Q(n584) );
  OR2X1 U597 ( .IN1(reg_b[20]), .IN2(n400), .Q(n518) );
  NAND2X0 U598 ( .IN1(n269), .IN2(n431), .QN(n223) );
  NOR2X0 U599 ( .IN1(reg_b[26]), .IN2(n419), .QN(n420) );
  NOR2X0 U600 ( .IN1(reg_b[24]), .IN2(n414), .QN(n415) );
  INVX0 U601 ( .IN(a_in[1]), .QN(n595) );
  INVX4 U602 ( .IN(n189), .QN(n237) );
  OA21X2 U603 ( .IN1(reg_a[1]), .IN2(n241), .IN3(n607), .Q(n226) );
  NOR2X0 U604 ( .IN1(reg_b[25]), .IN2(n417), .QN(n418) );
  NOR2X2 U605 ( .IN1(reg_b[15]), .IN2(n145), .QN(n232) );
  NBUFFX2 U606 ( .IN(n367), .Q(n342) );
  NBUFFX2 U607 ( .IN(reset_n), .Q(n367) );
  NBUFFX2 U608 ( .IN(reset_n), .Q(n366) );
  NBUFFX2 U609 ( .IN(reset_n), .Q(n365) );
  NBUFFX2 U610 ( .IN(reset_n), .Q(n364) );
  NBUFFX2 U611 ( .IN(reset_n), .Q(n363) );
  NBUFFX2 U612 ( .IN(reset_n), .Q(n362) );
  NBUFFX2 U613 ( .IN(reset_n), .Q(n361) );
  NBUFFX2 U614 ( .IN(reset_n), .Q(n360) );
  NBUFFX2 U615 ( .IN(reset_n), .Q(n359) );
  OR2X2 U616 ( .IN1(reg_b[9]), .IN2(n388), .Q(n450) );
  OA21X1 U617 ( .IN1(n469), .IN2(n468), .IN3(n467), .Q(n470) );
  AO222X1 U618 ( .IN1(n273), .IN2(reg_b[9]), .IN3(n182), .IN4(reg_a[9]), .IN5(
        b_in[9]), .IN6(n283), .Q(N101) );
  OA21X1 U619 ( .IN1(n577), .IN2(n209), .IN3(n576), .Q(n578) );
  NBUFFX2 U620 ( .IN(n186), .Q(n272) );
  AO222X1 U621 ( .IN1(n177), .IN2(reg_b[4]), .IN3(n182), .IN4(n103), .IN5(
        b_in[4]), .IN6(n277), .Q(N96) );
  AO22X1 U622 ( .IN1(n103), .IN2(n329), .IN3(result[4]), .IN4(n305), .Q(n93)
         );
  AO222X1 U623 ( .IN1(n275), .IN2(reg_b[2]), .IN3(n182), .IN4(n237), .IN5(
        b_in[2]), .IN6(n278), .Q(N94) );
  AO22X1 U624 ( .IN1(n237), .IN2(n330), .IN3(result[2]), .IN4(n306), .Q(n91)
         );
  MUX21X1 U625 ( .IN1(n550), .IN2(n549), .S(n557), .Q(n552) );
  NAND2X0 U626 ( .IN1(n160), .IN2(n579), .QN(n242) );
  NAND2X0 U627 ( .IN1(a_in[5]), .IN2(n109), .QN(n243) );
  NAND3X0 U628 ( .IN1(n242), .IN2(n243), .IN3(n134), .QN(N63) );
  NAND2X0 U629 ( .IN1(n160), .IN2(n441), .QN(n244) );
  NAND2X0 U630 ( .IN1(a_in[8]), .IN2(n108), .QN(n245) );
  NAND3X0 U631 ( .IN1(n244), .IN2(n245), .IN3(n128), .QN(N66) );
  NAND2X0 U632 ( .IN1(n160), .IN2(n514), .QN(n246) );
  NAND2X0 U633 ( .IN1(a_in[20]), .IN2(n191), .QN(n247) );
  NAND3X0 U634 ( .IN1(n246), .IN2(n247), .IN3(n127), .QN(N78) );
  OR4X1 U635 ( .IN1(reg_b[31]), .IN2(n179), .IN3(reg_b[4]), .IN4(reg_b[5]), 
        .Q(n59) );
  NAND2X0 U636 ( .IN1(n611), .IN2(n492), .QN(n248) );
  NAND2X0 U637 ( .IN1(a_in[17]), .IN2(n191), .QN(n249) );
  NAND3X0 U638 ( .IN1(n248), .IN2(n249), .IN3(n133), .QN(N75) );
  NAND2X0 U639 ( .IN1(n611), .IN2(n507), .QN(n250) );
  NAND2X0 U640 ( .IN1(a_in[19]), .IN2(n109), .QN(n251) );
  NAND3X0 U641 ( .IN1(n250), .IN2(n251), .IN3(n129), .QN(N77) );
  NAND2X0 U642 ( .IN1(n160), .IN2(n522), .QN(n252) );
  NAND3X0 U643 ( .IN1(n252), .IN2(n253), .IN3(n132), .QN(N79) );
  NAND2X0 U644 ( .IN1(n160), .IN2(n448), .QN(n254) );
  NAND2X0 U645 ( .IN1(a_in[9]), .IN2(n609), .QN(n255) );
  NAND3X0 U646 ( .IN1(n254), .IN2(n255), .IN3(n125), .QN(N67) );
  NAND2X0 U647 ( .IN1(reg_b[18]), .IN2(n391), .QN(n260) );
  AO222X1 U648 ( .IN1(n274), .IN2(reg_b[6]), .IN3(n182), .IN4(n236), .IN5(
        b_in[6]), .IN6(n277), .Q(N98) );
  OR4X1 U649 ( .IN1(reg_b[6]), .IN2(reg_b[7]), .IN3(reg_b[8]), .IN4(reg_b[9]), 
        .Q(n58) );
  OA21X1 U650 ( .IN1(n476), .IN2(n475), .IN3(n474), .Q(n477) );
  AO222X1 U651 ( .IN1(n177), .IN2(n258), .IN3(n182), .IN4(reg_a[11]), .IN5(
        b_in[11]), .IN6(n283), .Q(N103) );
  OA21X1 U652 ( .IN1(n483), .IN2(n482), .IN3(n481), .Q(n484) );
  NAND2X0 U653 ( .IN1(n160), .IN2(n585), .QN(n263) );
  NAND2X0 U654 ( .IN1(a_in[6]), .IN2(n609), .QN(n264) );
  NAND3X0 U655 ( .IN1(n263), .IN2(n264), .IN3(n131), .QN(N64) );
  NAND2X0 U656 ( .IN1(n160), .IN2(n528), .QN(n265) );
  NAND2X0 U657 ( .IN1(a_in[22]), .IN2(n108), .QN(n266) );
  NAND3X0 U658 ( .IN1(n265), .IN2(n266), .IN3(n130), .QN(N80) );
  AO22X1 U659 ( .IN1(n184), .IN2(n326), .IN3(result[1]), .IN4(n302), .Q(n98)
         );
  AO222X1 U660 ( .IN1(n275), .IN2(reg_b[28]), .IN3(n182), .IN4(reg_a[28]), 
        .IN5(b_in[28]), .IN6(n279), .Q(N120) );
  AO222X1 U661 ( .IN1(n273), .IN2(reg_b[24]), .IN3(n182), .IN4(reg_a[24]), 
        .IN5(b_in[24]), .IN6(n280), .Q(N116) );
  AO222X1 U662 ( .IN1(n274), .IN2(reg_b[15]), .IN3(n182), .IN4(reg_a[15]), 
        .IN5(b_in[15]), .IN6(n282), .Q(N107) );
  AO222X1 U663 ( .IN1(n273), .IN2(n179), .IN3(n182), .IN4(reg_a[3]), .IN5(
        b_in[3]), .IN6(n278), .Q(N95) );
  AO222X1 U664 ( .IN1(n274), .IN2(reg_b[10]), .IN3(n181), .IN4(reg_a[10]), 
        .IN5(b_in[10]), .IN6(n283), .Q(N102) );
  AO221X1 U665 ( .IN1(n611), .IN2(n610), .IN3(a_in[0]), .IN4(n609), .IN5(n608), 
        .Q(N58) );
  AO221X1 U666 ( .IN1(n611), .IN2(n587), .IN3(a_in[7]), .IN4(n108), .IN5(n586), 
        .Q(N65) );
  AO222X1 U667 ( .IN1(n272), .IN2(reg_b[22]), .IN3(n182), .IN4(reg_a[22]), 
        .IN5(b_in[22]), .IN6(n280), .Q(N114) );
  AO222X1 U668 ( .IN1(n274), .IN2(reg_b[7]), .IN3(n182), .IN4(n107), .IN5(
        b_in[7]), .IN6(n277), .Q(N99) );
  AO221X1 U669 ( .IN1(n160), .IN2(n486), .IN3(a_in[15]), .IN4(n108), .IN5(n485), .Q(N73) );
  AO22X1 U670 ( .IN1(n239), .IN2(reg_b[15]), .IN3(n165), .IN4(reg_a[15]), .Q(
        n485) );
  AO221X1 U671 ( .IN1(n611), .IN2(n546), .IN3(a_in[28]), .IN4(n191), .IN5(n545), .Q(N86) );
  AO22X1 U672 ( .IN1(n239), .IN2(reg_b[28]), .IN3(n165), .IN4(reg_a[28]), .Q(
        n545) );
  AO221X1 U673 ( .IN1(n611), .IN2(n540), .IN3(a_in[26]), .IN4(n108), .IN5(n539), .Q(N84) );
  AO22X1 U674 ( .IN1(n239), .IN2(reg_b[26]), .IN3(n165), .IN4(reg_a[26]), .Q(
        n539) );
  AO221X1 U675 ( .IN1(n160), .IN2(n534), .IN3(a_in[24]), .IN4(n191), .IN5(n533), .Q(N82) );
  AO22X1 U676 ( .IN1(n239), .IN2(reg_b[24]), .IN3(n165), .IN4(reg_a[24]), .Q(
        n533) );
  AO221X1 U677 ( .IN1(n611), .IN2(n500), .IN3(a_in[18]), .IN4(n609), .IN5(n499), .Q(N76) );
  AO22X1 U678 ( .IN1(n239), .IN2(reg_b[18]), .IN3(n166), .IN4(reg_a[18]), .Q(
        n499) );
  AO221X1 U679 ( .IN1(n611), .IN2(n479), .IN3(a_in[14]), .IN4(n109), .IN5(n478), .Q(N72) );
  AO22X1 U680 ( .IN1(n239), .IN2(reg_b[14]), .IN3(n166), .IN4(reg_a[14]), .Q(
        n478) );
  AO221X1 U681 ( .IN1(n160), .IN2(n458), .IN3(a_in[11]), .IN4(n609), .IN5(n457), .Q(N69) );
  AO22X1 U682 ( .IN1(n239), .IN2(n258), .IN3(n166), .IN4(reg_a[11]), .Q(n457)
         );
  AO221X1 U683 ( .IN1(n611), .IN2(n561), .IN3(a_in[30]), .IN4(n109), .IN5(n560), .Q(N88) );
  AO22X1 U684 ( .IN1(n239), .IN2(reg_b[30]), .IN3(n166), .IN4(reg_a[30]), .Q(
        n560) );
  AO221X1 U685 ( .IN1(n160), .IN2(n574), .IN3(a_in[4]), .IN4(n109), .IN5(n573), 
        .Q(N62) );
  AO22X1 U686 ( .IN1(n239), .IN2(reg_b[4]), .IN3(n166), .IN4(n103), .Q(n573)
         );
  AO221X1 U687 ( .IN1(n160), .IN2(n565), .IN3(a_in[2]), .IN4(n609), .IN5(n564), 
        .Q(N60) );
  AO22X1 U688 ( .IN1(n239), .IN2(reg_b[2]), .IN3(n165), .IN4(n237), .Q(n564)
         );
  AO221X1 U689 ( .IN1(n594), .IN2(n160), .IN3(a_in[31]), .IN4(n108), .IN5(n593), .Q(N89) );
  AO222X1 U690 ( .IN1(n275), .IN2(reg_b[1]), .IN3(n182), .IN4(n184), .IN5(
        b_in[1]), .IN6(n276), .Q(N93) );
  AO22X1 U691 ( .IN1(n239), .IN2(reg_b[7]), .IN3(n165), .IN4(n107), .Q(n586)
         );
  OA21X1 U692 ( .IN1(n505), .IN2(n504), .IN3(n503), .Q(n506) );
  INVX0 U693 ( .IN(n432), .QN(n269) );
  AO222X1 U694 ( .IN1(n177), .IN2(reg_b[31]), .IN3(n182), .IN4(reg_a[31]), 
        .IN5(b_in[31]), .IN6(n276), .Q(N123) );
  AO222X1 U695 ( .IN1(n273), .IN2(n262), .IN3(n182), .IN4(reg_a[16]), .IN5(
        b_in[16]), .IN6(n282), .Q(N108) );
  OA21X1 U696 ( .IN1(n512), .IN2(n511), .IN3(n510), .Q(n513) );
  OAI21X1 U697 ( .IN1(n520), .IN2(n519), .IN3(n518), .QN(n521) );
  AO22X1 U698 ( .IN1(n475), .IN2(n474), .IN3(reg_b[14]), .IN4(n370), .Q(n482)
         );
  AO221X1 U699 ( .IN1(n611), .IN2(n543), .IN3(a_in[27]), .IN4(n108), .IN5(n542), .Q(N85) );
  AO22X1 U700 ( .IN1(n239), .IN2(reg_b[27]), .IN3(n166), .IN4(reg_a[27]), .Q(
        n542) );
  AO221X1 U701 ( .IN1(n611), .IN2(n537), .IN3(a_in[25]), .IN4(n191), .IN5(n536), .Q(N83) );
  AO22X1 U702 ( .IN1(n239), .IN2(reg_b[25]), .IN3(n166), .IN4(reg_a[25]), .Q(
        n536) );
  AO221X1 U703 ( .IN1(n160), .IN2(n531), .IN3(a_in[23]), .IN4(n109), .IN5(n530), .Q(N81) );
  AO22X1 U704 ( .IN1(n239), .IN2(reg_b[23]), .IN3(n166), .IN4(reg_a[23]), .Q(
        n530) );
  AO221X1 U705 ( .IN1(n611), .IN2(n552), .IN3(a_in[29]), .IN4(n609), .IN5(n551), .Q(N87) );
  AO22X1 U706 ( .IN1(n239), .IN2(reg_b[29]), .IN3(n165), .IN4(reg_a[29]), .Q(
        n551) );
  AO221X1 U707 ( .IN1(n160), .IN2(n490), .IN3(a_in[16]), .IN4(n191), .IN5(n489), .Q(N74) );
  AO22X1 U708 ( .IN1(n239), .IN2(n262), .IN3(n166), .IN4(reg_a[16]), .Q(n489)
         );
  AO221X1 U709 ( .IN1(n611), .IN2(n464), .IN3(a_in[12]), .IN4(n109), .IN5(n463), .Q(N70) );
  AO22X1 U710 ( .IN1(n239), .IN2(n105), .IN3(n165), .IN4(n113), .Q(n463) );
  AO22X1 U711 ( .IN1(n504), .IN2(n503), .IN3(reg_b[19]), .IN4(n392), .Q(n511)
         );
  INVX4 U712 ( .IN(n439), .QN(n440) );
  AO221X1 U713 ( .IN1(n611), .IN2(n571), .IN3(a_in[3]), .IN4(n109), .IN5(n570), 
        .Q(N61) );
  AO22X1 U714 ( .IN1(n239), .IN2(n179), .IN3(n165), .IN4(reg_a[3]), .Q(n570)
         );
  AO221X1 U715 ( .IN1(n611), .IN2(n455), .IN3(a_in[10]), .IN4(n609), .IN5(n454), .Q(N68) );
  NBUFFX2 U716 ( .IN(n186), .Q(n275) );
  NBUFFX2 U717 ( .IN(n186), .Q(n274) );
  NBUFFX2 U718 ( .IN(n186), .Q(n273) );
  AND3X1 U719 ( .IN1(n114), .IN2(n338), .IN3(n588), .Q(gcd_ns[1]) );
  AO222X1 U720 ( .IN1(n273), .IN2(n176), .IN3(n182), .IN4(reg_a[0]), .IN5(
        b_in[0]), .IN6(n276), .Q(N92) );
  AO22X1 U721 ( .IN1(n239), .IN2(n176), .IN3(n166), .IN4(reg_a[0]), .Q(n608)
         );
  OR2X2 U722 ( .IN1(n439), .IN2(n111), .Q(n597) );
  NAND2X4 U723 ( .IN1(n390), .IN2(n389), .QN(n480) );
  NOR2X4 U724 ( .IN1(n487), .IN2(n205), .QN(n393) );
  NAND2X4 U725 ( .IN1(n399), .IN2(n398), .QN(n402) );
  NOR2X4 U726 ( .IN1(n402), .IN2(n401), .QN(n405) );
  NAND2X4 U727 ( .IN1(n523), .IN2(n403), .QN(n404) );
  NOR2X4 U728 ( .IN1(n405), .IN2(n404), .QN(n407) );
  NOR2X4 U729 ( .IN1(n407), .IN2(n406), .QN(n529) );
  NAND2X4 U730 ( .IN1(n408), .IN2(n409), .QN(n410) );
  NOR2X4 U731 ( .IN1(n158), .IN2(n420), .QN(n541) );
  NAND2X4 U732 ( .IN1(n421), .IN2(n422), .QN(n423) );
  OAI21X2 U733 ( .IN1(n433), .IN2(n284), .IN3(n434), .QN(n439) );
endmodule

